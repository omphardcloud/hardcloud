// hc_pkg.sv

package hc_pkg;
  import hc_user_pkg::*;

  // hardcloud internal definitions

  parameter HC_BUFFER_SIZE = HC_BUFFER_TX_SIZE + HC_BUFFER_RX_SIZE;

endpackage

