// hc_user_pkg.sv

package hc_user_pkg;

  //
  // HardCloud user definitions
  //

  parameter HC_BUFFER_TX_SIZE = 1;
  parameter HC_BUFFER_RX_SIZE = 1;

endpackage : hc_user_pkg

