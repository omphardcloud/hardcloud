// hc_user_pkg.sv

package hc_user_pkg;

  //
  // HardCloud user definitions
  //

  parameter HC_BUFFER_TX_SIZE = 1;
  parameter HC_BUFFER_RX_SIZE = 1;
  parameter HC_WRITE_FIFO_DEPTH = 1024;
  parameter HC_READ_REQUEST_FIFO_DEPTH = 8;

endpackage : hc_user_pkg

